package PE_pkg;

    typedef logic signed [15:0] int16_t;
    typedef logic signed [7:0] int8_t;

endpackage